/****************************************************
** RISC-V_B_instr.sv
** Author: Kai Roy, 
** Version: 1.0
** Date: 11/20/2023
** Description: This file handles the B Type instructions
** of a RISC-V Single Cycle Processor. (WIP)
****************************************************/
`timescale 1ns / 1ps
import riscv_pkg::*;

//Module for branch instructions
//- The new pc value is generated by this module
module B_type(
    input logic [31:0] instr,
	input logic [31:0] iaddr,
	input signed logic [31:0] imm,  rs1, rs2,
    output logic [31:0] pc
);
    import riscv_pkg::*;

	branch_instr branch;
    logic [31:0] u_rs1, u_rs2;

	assign u_rs1 = unsigned'(rs1);
	assign u_rs2 = unsigned'(rs2);
    assign branch = branch_instr'(instr[14:12])

    always_comb begin
		unique case(branch)
            BEQ:  out = (in1 == in2)     ? (iaddr+imm) : (iaddr+4);
            BNE:  out = (in1 != in2)     ? (iaddr+imm) : (iaddr+4);
            BLT:  out = (in1 < in2)      ? (iaddr+imm) : (iaddr+4);
            BGE:  out = (in1 >= in2)     ? (iaddr+imm) : (iaddr+4);
            BGEU: out = (u_rs1 < u_rs2)  ? (iaddr+imm) : (iaddr+4);
            BLTU: out = (u_rs1 >= u_rs2) ? (iaddr+imm) : (iaddr+4);
		endcase
	 end
endmodule