package rs_opcode; 
typedef enum logic [3:0] {rs0=4'b0000,rs1=4'b1000,rs2=4'b0001,rs3=4'b0010,rs4=4'b0011,rs5=4'b0100,rs6=4'b0101,rs7=4'b1101,rs8=4'b0110,rs9=4'b0111} OP_CODE_R;
endpackage